*T85T SPICE BSIM3 VERSION 3.1 PARAMETERS

*SPICE 3f5 Level 8, Star-HSPICE Level 49, UTMOST Level 8

* DATE: Sep  3/08
* LOT: T85T                  WAF: 2005
* Temperature_parameters=Default
.MODEL nm NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 3.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.485675
+K1      = 0.3634695      K2      = -0.0277136     K3      = 1E-3
+K3B     = 3.9409342      W0      = 1E-7           NLX     = 8.900764E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.2979753      DVT1    = 0.1605369      DVT2    = 0.2509178
+U0      = 436.2279588    UA      = -3.51975E-10   UB      = 3.216114E-18
+UC      = 4.919099E-10   VSAT    = 1.930256E5     A0      = 1.9922632
+AGS     = 0.7096599      B0      = 1.892162E-6    B1      = 5E-6
+KETA    = 0.05           A1      = 7.799989E-4    A2      = 0.3
+RDSW    = 150            PRWG    = 0.3506787      PRWB    = 0.1097886
+WR      = 1              WINT    = 7.71429E-9     LINT    = 1.039368E-8
+DWG     = 1.205322E-8    DWB     = 8.815731E-9    VOFF    = -0.0331648
+NFACTOR = 2.5            CIT     = 0              CDSC    = 2.4E-4
+CDSCD   = 0              CDSCB   = 0              ETA0    = 2.754257E-6
+ETAB    = -0.0108095     DSUB    = 4.0643E-6      PCLM    = 1.9769478
+PDIBLC1 = 0.9710894      PDIBLC2 = 0.01           PDIBLCB = 0.1
+DROUT   = 0.9993653      PSCBE1  = 7.973288E10    PSCBE2  = 5.02618E-10
+PVAG    = 0.536394       DELTA   = 0.01           RSH     = 6.7
+MOBMOD  = 1              PRT     = 0              UTE     = -1.5
+KT1     = -0.11          KT1L    = 0              KT2     = 0.022
+UA1     = 4.31E-9        UB1     = -7.61E-18      UC1     = -5.6E-11
+AT      = 3.3E4          WL      = 0              WLN     = 1
+WW      = 0              WWN     = 1              WWL     = 0
+LL      = 0              LLN     = 1              LW      = 0
+LWN     = 1              LWL     = 0              CAPMOD  = 2
+XPART   = 0.5            CGDO    = 3.74E-10       CGSO    = 3.74E-10
+CGBO    = 1E-12          CJ      = 9.581316E-4    PB      = 0.9759771
+MJ      = 0.404514       CJSW    = 1E-10          PBSW    = 0.8002028
+MJSW    = 0.6            CJSWG   = 3.3E-10        PBSWG   = 0.8002028
+MJSWG   = 0.6            CF      = 0              PVTH0   = 2.009264E-4
+PRDSW   = 0              PK2     = 1.30501E-3     WKETA   = 7.565815E-3
+LKETA   = 0.0327047      PU0     = 4.4729531      PUA     = 1.66833E-11
+PUB     = 0              PVSAT   = 653.2294237    PETA0   = 1E-4
+PKETA   = -0.0101124      )
*
.MODEL pm PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 3.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.2156906
+K1      = 0.2680989      K2      = 4.539197E-3    K3      = 0.097375
+K3B     = 6.5043674      W0      = 1E-6           NLX     = 2.836757E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0              DVT1    = 1              DVT2    = 0.1
+U0      = 106.670318     UA      = 1.152986E-9    UB      = 2.377339E-21
+UC      = -1.93766E-11   VSAT    = 1.190739E5     A0      = 1.7356069
+AGS     = 0.6166218      B0      = 7.467707E-6    B1      = 4.992767E-6
+KETA    = 0.0157125      A1      = 8.723417E-3    A2      = 0.8713799
+RDSW    = 105            PRWG    = -0.5           PRWB    = 0.5
+WR      = 1              WINT    = 0              LINT    = 1.495916E-8
+DWG     = 6.058254E-9    DWB     = -1.83713E-8    VOFF    = -0.1022829
+NFACTOR = 1.5332272      CIT     = 0              CDSC    = 2.4E-4
+CDSCD   = 0              CDSCB   = 0              ETA0    = 0.0110506
+ETAB    = -2.941775E-3   DSUB    = 2.419246E-3    PCLM    = 0.2085802
+PDIBLC1 = 9.972716E-4    PDIBLC2 = -1.39497E-13   PDIBLCB = -1E-3
+DROUT   = 0.6860806      PSCBE1  = 1.849353E9     PSCBE2  = 5.675435E-10
+PVAG    = 0.0149584      DELTA   = 0.01           RSH     = 6.6
+MOBMOD  = 1              PRT     = 0              UTE     = -1.5
+KT1     = -0.11          KT1L    = 0              KT2     = 0.022
+UA1     = 4.31E-9        UB1     = -7.61E-18      UC1     = -5.6E-11
+AT      = 3.3E4          WL      = 0              WLN     = 1
+WW      = 0              WWN     = 1              WWL     = 0
+LL      = 0              LLN     = 1              LW      = 0
+LWN     = 1              LWL     = 0              CAPMOD  = 2
+XPART   = 0.5            CGDO    = 3.42E-10       CGSO    = 3.42E-10
+CGBO    = 1E-12          CJ      = 1.15643E-3     PB      = 0.8
+MJ      = 0.4399866      CJSW    = 1.133806E-10   PBSW    = 0.8
+MJSW    = 0.1146401      CJSWG   = 4.22E-10       PBSWG   = 0.8
+MJSWG   = 0.1146401      CF      = 0              PVTH0   = 1.282832E-3
+PRDSW   = 44.1361752     PK2     = 2.459655E-3    WKETA   = 0.0352131
+LKETA   = 0.0128331      PU0     = -1.2608844     PUA     = -4.27994E-11
+PUB     = 1.628153E-28   PVSAT   = -50            PETA0   = 7.039749E-5
+PKETA   = -5.052402E-3    )
