* 741 OPAMP Testbench
* Hisham Elreedy
*----------------------------------------------------
*	Models and Parameters
*----------------------------------------------------
.include 'LM741.MOD'

*---------------------------------------------------
*	Netlist, Circuit Elements and Signal Sources
*---------------------------------------------------
V1 v1 gnd 1V


*--------------------------------------------------
*	Stimulus and Simulation
*--------------------------------------------------
.op

.end
